module top_module( input in, output out );
    // assign (output) = (input)
    assign out = in;

endmodule